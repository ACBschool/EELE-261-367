library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity top is 

	port(SW 		: in std_logic_vector(7 downto 0);
		  LEDR	: out std_logic_vector(9 downto 0);
		  HEX0	: out std_logic_vector(6 downto 0);
		  HEX1 	: out std_logic_vector(6 downto 0);
		  HEX2	: out std_logic_vector(6 downto 0);
		  HEX3	: out std_logic_vector(6 downto 0);
		  HEX4	: out std_logic_vector(6 downto 0);
		  HEX5 	: out std_logic_vector(6 downto 0));

end entity;


architecture top_arch of top is


------------------------------------------------------------------------------------------------
-------------------------------Component-Subsystems---------------------------------------------
------------------------------------------------------------------------------------------------

	-- hex decoder component
	component char_decoder
		port(BIN_IN		: in std_logic_vector (3 downto 0);
			  HEX_OUT	: out std_logic_vector ( 6 downto 0));
	end component;
	
	


	
	
------------------------------------------------------------------------------------------------	
---------------------------Internal-signals-----------------------------------------------------
------------------------------------------------------------------------------------------------

	signal Carry : std_logic;	--interim signal to hold the carry bit. Descriptive.a
	signal Sum	 : std_logic_vector(3 downto 0);	-- interim hold sum of adder.
	signal Sum_uns : unsigned(4 downto 0);
	
	
------------------------------------------------------------------------------------------------	
------------------------------------------------------------------------------------------------
-------------------Begin-Modeling---------------------------------------------------------------
------------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------------


	
	begin

	
------------------------------------------------------------------------------------------------
------------------------------------------General-Assignment-I/O--------------------------------
------------------------------------------------------------------------------------------------

		LEDR(7 downto 0) <= SW;
		LEDR(9) <= Carry;

------------------------------------------------------------------------------------------------
--------------------------------------HEX-displays-subsystem------------------------------------
------------------------------------------------------------------------------------------------

	-- HEX component instantiation
	
		C0	: char_decoder port map ( BIN_IN => SW(3 downto 0) , HEX_OUT => HEX0);
		C2	: char_decoder port map ( BIN_IN => SW(7 downto 4) , HEX_OUT => HEX2);
		HEX1 <= "1111111";
		HEX3 <= "1111111";
		C4	: char_decoder port map ( BIN_IN => Sum(3 downto 0) , HEX_OUT => HEX4);
		C5	: char_decoder port map ( BIN_IN => "000" & Carry , HEX_OUT => HEX5);



------------------------------------------------------------------------------------------------
-------------------------------Adder-Subsystem--------------------------------------------------
------------------------------------------------------------------------------------------------

		Sum_uns <= unsigned(('0' & SW(7 downto 4))) + unsigned(('0' & SW(3 downto 0)));

		Sum <= std_logic_vector(Sum_uns(3 downto 0));
		Carry <= Sum_uns(4);


------------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------------


end architecture;
	




