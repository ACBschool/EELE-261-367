library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom_4x4_async is
	port (address	: in std_logic_vector(1 downto 0);
	      clock	: in std_logic;
	      data_out	: out std_logic_vector(3 downto 0));
end entity;


architecture rom_4x4_async_arch of rom_4x4_async is

			--   array indices, what is contained with each index
	type ROM_type is array (0 to 3) of std_logic_vector(3 downto 0);

	constant ROM : ROM_type := (0 => "1110", -- read as address zero contains 1110
			      1 => "0010",
			      2 => "1111",
			      3 => "0100");
	begin


	--data_out <= ROM(to_integer(unsigned(address))); just this if asynchronous

	SYNC_PROC : process(clock)	-- process of synchronous update
		begin
			if(rising_edge(clock)) then
				data_out <= ROM(to_integer(unsigned(address)));	
			end if;
	end process;

end architecture;
